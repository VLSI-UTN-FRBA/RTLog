module fir_transpose
	(
		input wire rst,
		input wire clk,
		input wire [15:0] X,
		output reg [15:0] Y,
	);

	wire net_tie_hi;
	wire net_ti_lo;
	reg q_19;
	reg q_21;
	reg q_23;
	reg q_25;
	reg q_27;
	reg q_29;
	reg q_31;
	reg q_33;
	reg q_35;
	reg q_37;
	reg q_39;
	reg q_41;
	reg q_43;
	reg q_45;
	reg q_47;
	reg q_49;
	wire buf_50;
	wire buf_51;
	wire buf_52;
	wire buf_53;
	wire buf_54;
	wire buf_55;
	wire buf_56;
	wire buf_57;
	wire buf_58;
	wire buf_59;
	wire buf_60;
	wire buf_61;
	wire buf_62;
	wire buf_63;
	wire buf_64;
	wire buf_65;
	wire buf_66;
	wire buf_67;
	wire buf_68;
	wire buf_69;
	wire buf_70;
	wire buf_71;
	wire buf_72;
	wire buf_73;
	wire buf_74;
	wire buf_75;
	wire buf_76;
	wire buf_77;
	wire buf_78;
	wire buf_79;
	wire buf_80;
	wire buf_81;
	wire buf_82;
	wire buf_83;
	wire buf_84;
	wire buf_85;
	wire buf_86;
	wire buf_87;
	wire buf_88;
	wire buf_89;
	wire buf_90;
	wire buf_91;
	wire buf_92;
	wire buf_93;
	wire buf_94;
	wire buf_95;
	wire buf_96;
	wire buf_97;
	wire buf_98;
	wire buf_99;
	wire buf_100;
	wire buf_101;
	wire buf_102;
	wire buf_103;
	wire buf_104;
	wire buf_105;
	wire buf_106;
	wire buf_107;
	wire buf_108;
	wire buf_109;
	wire buf_110;
	wire buf_111;
	wire buf_112;
	wire buf_113;
	wire buf_114;
	wire buf_115;
	wire buf_116;
	wire buf_117;
	wire buf_118;
	wire buf_119;
	wire buf_120;
	wire buf_121;
	wire buf_122;
	wire buf_123;
	wire buf_124;
	wire buf_125;
	wire buf_126;
	wire buf_127;
	wire buf_128;
	wire buf_129;
	wire buf_130;
	wire buf_131;
	wire buf_132;
	wire buf_133;
	wire buf_134;
	wire buf_135;
	wire buf_136;
	wire buf_137;
	wire buf_138;
	wire buf_139;
	wire buf_140;
	wire buf_141;
	wire buf_142;
	wire buf_143;
	wire buf_144;
	wire buf_145;
	wire buf_146;
	wire buf_147;
	wire buf_148;
	wire buf_149;
	wire buf_150;
	wire buf_151;
	wire buf_152;
	wire buf_153;
	wire buf_154;
	wire buf_155;
	wire buf_156;
	wire buf_157;
	wire buf_158;
	wire buf_159;
	wire buf_160;
	wire buf_161;
	wire buf_162;
	wire buf_163;
	wire buf_164;
	wire buf_165;
	wire buf_166;
	wire buf_167;
	wire buf_168;
	wire buf_169;
	wire buf_170;
	wire buf_171;
	wire buf_172;
	wire buf_173;
	wire buf_174;
	wire buf_175;
	wire buf_176;
	wire buf_177;
	wire buf_178;
	wire buf_179;
	wire buf_180;
	wire buf_181;
	wire buf_182;
	wire buf_183;
	wire buf_184;
	wire buf_185;
	wire buf_186;
	wire buf_187;
	wire buf_188;
	wire buf_189;
	wire buf_190;
	wire buf_191;
	wire buf_192;
	wire buf_193;
	wire buf_194;
	wire buf_195;
	wire buf_196;
	wire buf_197;
	wire buf_198;
	wire buf_199;
	wire buf_200;
	wire buf_201;
	wire buf_202;
	wire buf_203;
	wire buf_204;
	wire buf_205;
	wire buf_206;
	wire buf_207;
	wire buf_208;
	wire buf_209;
	wire buf_210;
	wire buf_211;
	wire buf_212;
	wire buf_213;
	wire buf_214;
	wire buf_215;
	wire buf_216;
	wire buf_217;
	wire buf_218;
	wire buf_219;
	wire buf_220;
	wire buf_221;
	wire buf_222;
	wire buf_223;
	wire buf_224;
	wire buf_225;
	wire buf_226;
	wire buf_227;
	wire buf_228;
	wire buf_229;
	wire buf_230;
	wire buf_231;
	wire buf_232;
	wire buf_233;
	wire buf_234;
	wire buf_235;
	wire buf_236;
	wire buf_237;
	wire buf_238;
	wire buf_239;
	wire buf_240;
	wire buf_241;
	wire buf_242;
	wire buf_243;
	wire buf_244;
	wire buf_245;
	wire buf_246;
	wire buf_247;
	wire buf_248;
	wire buf_249;
	wire buf_250;
	wire buf_251;
	wire buf_252;
	wire buf_253;
	wire buf_254;
	wire buf_255;
	wire buf_256;
	wire buf_257;
	wire buf_258;
	wire buf_259;
	wire buf_260;
	wire buf_261;
	wire buf_262;
	wire buf_263;
	wire buf_264;
	wire buf_265;
	wire buf_266;
	wire buf_267;
	wire buf_268;
	wire buf_269;
	wire buf_270;
	wire buf_271;
	wire buf_272;
	wire buf_273;
	wire buf_274;
	wire buf_275;
	wire buf_276;
	wire buf_277;
	wire buf_278;
	wire buf_279;
	wire buf_280;
	wire buf_281;
	wire buf_282;
	wire buf_283;
	wire buf_284;
	wire buf_285;
	wire buf_286;
	wire buf_287;
	wire buf_288;
	wire buf_289;
	reg q_290;
	reg q_291;
	reg q_292;
	reg q_293;
	reg q_294;
	reg q_295;
	reg q_296;
	reg q_297;
	reg q_298;
	reg q_299;
	reg q_300;
	reg q_301;
	reg q_302;
	reg q_303;
	reg q_304;
	reg q_305;
	reg q_306;
	reg q_307;
	reg q_308;
	reg q_309;
	reg q_310;
	reg q_311;
	reg q_312;
	reg q_313;
	reg q_314;
	reg q_315;
	reg q_316;
	reg q_317;
	reg q_318;
	reg q_319;
	reg q_320;
	reg q_321;
	reg q_322;
	reg q_323;
	reg q_324;
	reg q_325;
	reg q_326;
	reg q_327;
	reg q_328;
	reg q_329;
	reg q_330;
	reg q_331;
	reg q_332;
	reg q_333;
	reg q_334;
	reg q_335;
	reg q_336;
	reg q_337;
	reg q_338;
	reg q_339;
	reg q_340;
	reg q_341;
	reg q_342;
	reg q_343;
	reg q_344;
	reg q_345;
	reg q_346;
	reg q_347;
	reg q_348;
	reg q_349;
	reg q_350;
	reg q_351;
	reg q_352;
	reg q_353;
	wire mult_354[31:0];
	wire mult_355[31:0];
	wire mult_356[31:0];
	wire mult_357[31:0];
	wire add_358[15:0];
	wire add_359[15:0];
	wire add_360[15:0];
	wire net_0;
	wire net_1;
	wire net_2;
	wire net_3;
	wire net_4;
	wire net_5;
	wire net_6;
	wire net_7;
	wire net_8;
	wire net_9;
	wire net_10;
	wire net_11;
	wire net_12;
	wire net_13;
	wire net_14;
	wire net_15;
	wire net_16;
	wire net_17;
	wire net_18;
	wire net_19;
	wire net_20;
	wire net_21;
	wire net_22;
	wire net_23;
	wire net_24;
	wire net_25;
	wire net_26;
	wire net_27;
	wire net_28;
	wire net_29;
	wire net_30;
	wire net_31;
	wire net_32;
	wire net_33;
	wire net_34;
	wire net_35;
	wire net_36;
	wire net_37;
	wire net_38;
	wire net_39;
	wire net_40;
	wire net_41;
	wire net_42;
	wire net_43;
	wire net_44;
	wire net_45;
	wire net_46;
	wire net_47;
	wire net_48;
	wire net_49;
	wire net_50;
	wire net_51;
	wire net_52;
	wire net_53;
	wire net_54;
	wire net_55;
	wire net_56;
	wire net_57;
	wire net_58;
	wire net_59;
	wire net_60;
	wire net_61;
	wire net_62;
	wire net_63;
	wire net_64;
	wire net_65;
	wire net_66;
	wire net_67;
	wire net_68;
	wire net_69;
	wire net_70;
	wire net_71;
	wire net_72;
	wire net_73;
	wire net_74;
	wire net_75;
	wire net_76;
	wire net_77;
	wire net_78;
	wire net_79;
	wire net_80;
	wire net_81;
	wire net_82;
	wire net_83;
	wire net_84;
	wire net_85;
	wire net_86;
	wire net_87;
	wire net_88;
	wire net_89;
	wire net_90;
	wire net_91;
	wire net_92;
	wire net_93;
	wire net_94;
	wire net_95;
	wire net_96;
	wire net_97;
	wire net_98;
	wire net_99;
	wire net_100;
	wire net_101;
	wire net_102;
	wire net_103;
	wire net_104;
	wire net_105;
	wire net_106;
	wire net_107;
	wire net_108;
	wire net_109;
	wire net_110;
	wire net_111;
	wire net_112;
	wire net_113;
	wire net_114;
	wire net_115;
	wire net_116;
	wire net_117;
	wire net_118;
	wire net_119;
	wire net_120;
	wire net_121;
	wire net_122;
	wire net_123;
	wire net_124;
	wire net_125;
	wire net_126;
	wire net_127;
	wire net_128;
	wire net_129;
	wire net_130;
	wire net_131;
	wire net_132;
	wire net_133;
	wire net_134;
	wire net_135;
	wire net_136;
	wire net_137;
	wire net_138;
	wire net_139;
	wire net_140;
	wire net_141;
	wire net_142;
	wire net_143;
	wire net_144;
	wire net_145;
	wire net_146;
	wire net_147;
	wire net_148;
	wire net_149;
	wire net_150;
	wire net_151;
	wire net_152;
	wire net_153;
	wire net_154;
	wire net_155;
	wire net_156;
	wire net_157;
	wire net_158;
	wire net_159;
	wire net_160;
	wire net_161;
	wire net_162;
	wire net_163;
	wire net_164;
	wire net_165;
	wire net_166;
	wire net_167;
	wire net_168;
	wire net_169;
	wire net_170;
	wire net_171;
	wire net_172;
	wire net_173;
	wire net_174;
	wire net_175;
	wire net_176;
	wire net_177;
	wire net_178;
	wire net_179;
	wire net_180;
	wire net_181;
	wire net_182;
	wire net_183;
	wire net_184;
	wire net_185;
	wire net_186;
	wire net_187;
	wire net_188;
	wire net_189;
	wire net_190;
	wire net_191;
	wire net_192;
	wire net_193;
	wire net_194;
	wire net_195;
	wire net_196;
	wire net_197;
	wire net_198;
	wire net_199;
	wire net_200;
	wire net_201;
	wire net_202;
	wire net_203;
	wire net_204;
	wire net_205;
	wire net_206;
	wire net_207;
	wire net_208;
	wire net_209;
	wire net_210;
	wire net_211;
	wire net_212;
	wire net_213;
	wire net_214;
	wire net_215;
	wire net_216;
	wire net_217;
	wire net_218;
	wire net_219;
	wire net_220;
	wire net_221;
	wire net_222;
	wire net_223;
	wire net_224;
	wire net_225;
	wire net_226;
	wire net_227;
	wire net_228;
	wire net_229;
	wire net_230;
	wire net_231;
	wire net_232;
	wire net_233;
	wire net_234;
	wire net_235;
	wire net_236;
	wire net_237;
	wire net_238;
	wire net_239;
	wire net_240;
	wire net_241;
	wire net_242;
	wire net_243;
	wire net_244;
	wire net_245;
	wire net_246;
	wire net_247;
	wire net_248;
	wire net_249;
	wire net_250;
	wire net_251;
	wire net_252;
	wire net_253;
	wire net_254;
	wire net_255;
	wire net_256;
	wire net_257;
	wire net_258;
	wire net_259;
	wire net_260;
	wire net_261;
	wire net_262;
	wire net_263;
	wire net_264;
	wire net_265;
	wire net_266;
	wire net_267;
	wire net_268;
	wire net_269;
	wire net_270;
	wire net_271;
	wire net_272;
	wire net_273;
	wire net_274;
	wire net_275;
	wire net_276;
	wire net_277;
	wire net_278;
	wire net_279;
	wire net_280;
	wire net_281;
	wire net_282;
	wire net_283;
	wire net_284;
	wire net_285;
	wire net_286;
	wire net_287;
	wire net_288;
	wire net_289;
	wire net_290;
	wire net_291;
	wire net_292;
	wire net_293;
	wire net_294;
	wire net_295;
	wire net_296;
	wire net_297;
	wire net_298;
	wire net_299;
	wire net_300;
	wire net_301;
	wire net_302;
	wire net_303;
	wire net_304;
	wire net_305;
	wire net_306;
	wire net_307;
	wire net_308;
	wire net_309;
	wire net_310;
	wire net_311;
	wire net_312;
	wire net_313;
	wire net_314;
	wire net_315;
	wire net_316;
	wire net_317;
	wire net_318;
	wire net_319;
	wire net_320;
	wire net_321;
	wire net_322;
	wire net_323;
	wire net_324;
	wire net_325;
	wire net_326;
	wire net_327;
	wire net_328;
	wire net_329;
	wire net_330;
	wire net_331;
	wire net_332;
	wire net_333;
	wire net_334;
	wire net_335;
	wire net_336;
	wire net_337;
	wire net_338;
	wire net_339;
	wire net_340;
	wire net_341;
	wire net_342;
	wire net_343;
	wire net_344;
	wire net_345;
	wire net_346;
	wire net_347;
	wire net_348;
	wire net_349;
	wire net_350;
	wire net_351;
	wire net_352;
	wire net_353;
	wire net_354;
	wire net_355;
	wire net_356;
	wire net_357;
	wire net_358;
	wire net_359;
	wire net_360;
	wire net_361;
	wire net_362;
	wire net_363;
	wire net_364;
	wire net_365;
	wire net_366;
	wire net_367;
	wire net_368;
	wire net_369;
	wire net_370;
	wire net_371;
	wire net_372;
	wire net_373;
	wire net_374;
	wire net_375;
	wire net_376;
	wire net_377;
	wire net_378;
	wire net_379;
	wire net_380;
	wire net_381;
	wire net_382;
	wire net_383;
	wire net_384;
	wire net_385;
	wire net_386;
	wire net_387;
	wire net_388;
	wire net_389;
	wire net_390;
	wire net_391;
	wire net_392;
	wire net_393;
	wire net_394;
	wire net_395;
	wire net_396;
	wire net_397;
	wire net_398;
	wire net_399;
	wire net_400;
	wire net_401;
	wire net_402;
	wire net_403;
	wire net_404;
	wire net_405;
	wire net_406;
	wire net_407;
	wire net_408;
	wire net_409;
	wire net_410;
	wire net_411;
	wire net_412;
	wire net_413;
	wire net_414;
	wire net_415;
	wire net_416;
	wire net_417;
	wire net_418;
	wire net_419;
	wire net_420;
	wire net_421;
	wire net_422;
	wire net_423;
	wire net_424;
	wire net_425;
	wire net_426;
	wire net_427;
	wire net_428;
	wire net_429;
	wire net_430;
	wire net_431;
	wire net_432;
	wire net_433;
	wire net_434;
	wire net_435;
	wire net_436;
	wire net_437;
	wire net_438;
	wire net_439;
	wire net_440;
	wire net_441;
	wire net_442;
	wire net_443;
	wire net_444;
	wire net_445;
	wire net_446;
	wire net_447;
	wire net_448;
	wire net_449;
	wire net_450;
	wire net_451;
	wire net_452;
	wire net_453;
	wire net_454;
	wire net_455;
	wire net_456;
	wire net_457;
	wire net_458;
	wire net_459;
	wire net_460;
	wire net_461;
	wire net_462;
	wire net_463;
	wire net_464;
	wire net_465;
	wire net_466;
	wire net_467;
	wire net_468;
	wire net_469;
	wire net_470;
	wire net_471;
	wire net_472;
	wire net_473;
	wire net_474;
	wire net_475;
	wire net_476;
	wire net_477;
	wire net_478;
	wire net_479;
	wire net_480;
	wire net_481;
	wire net_482;
	wire net_483;
	wire net_484;
	wire net_485;
	wire net_486;
	wire net_487;
	wire net_488;
	wire net_489;
	wire net_490;
	wire net_491;
	wire net_492;
	wire net_493;
	wire net_494;
	wire net_495;
	wire net_496;
	wire net_497;
	wire net_498;
	wire net_499;
	wire net_500;
	wire net_501;
	wire net_502;
	wire net_503;
	wire net_504;
	wire net_505;
	wire net_506;
	wire net_507;
	wire net_508;
	wire net_509;
	wire net_510;
	wire net_511;
	wire net_512;
	wire net_513;
	wire net_514;
	wire net_515;
	wire net_516;
	wire net_517;
	wire net_518;
	wire net_519;
	wire net_520;
	wire net_521;
	wire net_522;
	wire net_523;
	wire net_524;
	wire net_525;
	wire net_526;
	wire net_527;
	wire net_528;
	wire net_529;
	wire net_530;
	wire net_531;
	wire net_532;
	wire net_533;
	wire net_534;
	wire net_535;
	wire net_536;
	wire net_537;
	wire net_538;
	wire net_539;
	wire net_540;
	wire net_541;
	wire net_542;
	wire net_543;
	wire net_544;
	wire net_545;
	wire net_546;
	wire net_547;
	wire net_548;
	wire net_549;
	wire net_550;
	wire net_551;
	wire net_552;
	wire net_553;
	wire net_554;
	wire net_555;
	wire net_556;
	wire net_557;
	wire net_558;
	wire net_559;

	assign net_tie_hi = 1'b1;
	assign net_ti_lo = 1'b0;
	assign net_16 = net_tie_lo;
	assign net_18 = net_tie_lo;
	assign net_29 = net_tie_lo;
	assign net_30 = net_tie_lo;
	assign net_31 = net_tie_lo;
	assign net_32 = net_tie_lo;
	assign net_34 = net_tie_lo;
	assign net_45 = net_tie_lo;
	assign net_46 = net_tie_lo;
	assign net_47 = net_tie_lo;
	assign net_49 = net_tie_lo;
	assign net_53 = net_tie_lo;
	assign net_54 = net_tie_lo;
	assign net_57 = net_tie_lo;
	assign net_58 = net_tie_lo;
	assign net_59 = net_tie_lo;
	assign net_60 = net_tie_lo;
	assign net_61 = net_tie_lo;
	assign net_62 = net_tie_lo;
	assign net_63 = net_tie_lo;
	assign net_64 = net_tie_lo;
	assign net_66 = net_tie_lo;
	assign net_77 = net_tie_lo;
	assign net_78 = net_tie_lo;
	assign net_79 = net_tie_lo;
	assign net_17 = net_tie_hi;
	assign net_19 = net_tie_hi;
	assign net_20 = net_tie_hi;
	assign net_21 = net_tie_hi;
	assign net_22 = net_tie_hi;
	assign net_23 = net_tie_hi;
	assign net_24 = net_tie_hi;
	assign net_25 = net_tie_hi;
	assign net_26 = net_tie_hi;
	assign net_27 = net_tie_hi;
	assign net_28 = net_tie_hi;
	assign net_33 = net_tie_hi;
	assign net_35 = net_tie_hi;
	assign net_36 = net_tie_hi;
	assign net_37 = net_tie_hi;
	assign net_38 = net_tie_hi;
	assign net_39 = net_tie_hi;
	assign net_40 = net_tie_hi;
	assign net_41 = net_tie_hi;
	assign net_42 = net_tie_hi;
	assign net_43 = net_tie_hi;
	assign net_44 = net_tie_hi;
	assign net_48 = net_tie_hi;
	assign net_50 = net_tie_hi;
	assign net_51 = net_tie_hi;
	assign net_52 = net_tie_hi;
	assign net_55 = net_tie_hi;
	assign net_56 = net_tie_hi;
	assign net_65 = net_tie_hi;
	assign net_67 = net_tie_hi;
	assign net_68 = net_tie_hi;
	assign net_69 = net_tie_hi;
	assign net_70 = net_tie_hi;
	assign net_71 = net_tie_hi;
	assign net_72 = net_tie_hi;
	assign net_73 = net_tie_hi;
	assign net_74 = net_tie_hi;
	assign net_75 = net_tie_hi;
	assign net_76 = net_tie_hi;
	assign net_80 = X[0];
	assign net_81 = X[1];
	assign net_82 = X[2];
	assign net_83 = X[3];
	assign net_84 = X[4];
	assign net_85 = X[5];
	assign net_86 = X[6];
	assign net_87 = X[7];
	assign net_88 = X[8];
	assign net_89 = X[9];
	assign net_90 = X[10];
	assign net_91 = X[11];
	assign net_92 = X[12];
	assign net_93 = X[13];
	assign net_94 = X[14];
	assign net_95 = X[15];
	assign Y[0] = net_0;
	assign net_0 = q_19;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_19 = 1'b0;
		end
		else
		begin
			q_19 = net_544;
		end
	end

	assign Y[1] = net_1;
	assign net_1 = q_21;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_21 = 1'b0;
		end
		else
		begin
			q_21 = net_545;
		end
	end

	assign Y[2] = net_2;
	assign net_2 = q_23;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_23 = 1'b0;
		end
		else
		begin
			q_23 = net_546;
		end
	end

	assign Y[3] = net_3;
	assign net_3 = q_25;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_25 = 1'b0;
		end
		else
		begin
			q_25 = net_547;
		end
	end

	assign Y[4] = net_4;
	assign net_4 = q_27;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_27 = 1'b0;
		end
		else
		begin
			q_27 = net_548;
		end
	end

	assign Y[5] = net_5;
	assign net_5 = q_29;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_29 = 1'b0;
		end
		else
		begin
			q_29 = net_549;
		end
	end

	assign Y[6] = net_6;
	assign net_6 = q_31;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_31 = 1'b0;
		end
		else
		begin
			q_31 = net_550;
		end
	end

	assign Y[7] = net_7;
	assign net_7 = q_33;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_33 = 1'b0;
		end
		else
		begin
			q_33 = net_551;
		end
	end

	assign Y[8] = net_8;
	assign net_8 = q_35;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_35 = 1'b0;
		end
		else
		begin
			q_35 = net_552;
		end
	end

	assign Y[9] = net_9;
	assign net_9 = q_37;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_37 = 1'b0;
		end
		else
		begin
			q_37 = net_553;
		end
	end

	assign Y[10] = net_10;
	assign net_10 = q_39;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_39 = 1'b0;
		end
		else
		begin
			q_39 = net_554;
		end
	end

	assign Y[11] = net_11;
	assign net_11 = q_41;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_41 = 1'b0;
		end
		else
		begin
			q_41 = net_555;
		end
	end

	assign Y[12] = net_12;
	assign net_12 = q_43;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_43 = 1'b0;
		end
		else
		begin
			q_43 = net_556;
		end
	end

	assign Y[13] = net_13;
	assign net_13 = q_45;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_45 = 1'b0;
		end
		else
		begin
			q_45 = net_557;
		end
	end

	assign Y[14] = net_14;
	assign net_14 = q_47;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_47 = 1'b0;
		end
		else
		begin
			q_47 = net_558;
		end
	end

	assign Y[15] = net_15;
	assign net_15 = q_49;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_49 = 1'b0;
		end
		else
		begin
			q_49 = net_559;
		end
	end


	assign buf_50 = net_320;


	assign buf_51 = net_321;


	assign buf_52 = net_322;


	assign buf_53 = net_323;


	assign buf_54 = net_324;


	assign buf_55 = net_325;


	assign buf_56 = net_326;


	assign buf_57 = net_327;


	assign buf_58 = net_328;


	assign buf_59 = net_329;


	assign buf_60 = net_330;


	assign buf_61 = net_331;


	assign buf_62 = net_332;


	assign buf_63 = net_333;


	assign buf_64 = net_334;


	assign buf_65 = net_335;

	assign net_352 = buf_66;

	assign buf_66 = net_336;

	assign net_353 = buf_67;

	assign buf_67 = net_337;

	assign net_354 = buf_68;

	assign buf_68 = net_338;

	assign net_355 = buf_69;

	assign buf_69 = net_339;

	assign net_356 = buf_70;

	assign buf_70 = net_340;

	assign net_357 = buf_71;

	assign buf_71 = net_341;

	assign net_358 = buf_72;

	assign buf_72 = net_342;

	assign net_359 = buf_73;

	assign buf_73 = net_343;

	assign net_360 = buf_74;

	assign buf_74 = net_344;

	assign net_361 = buf_75;

	assign buf_75 = net_345;

	assign net_362 = buf_76;

	assign buf_76 = net_346;

	assign net_363 = buf_77;

	assign buf_77 = net_347;

	assign net_364 = buf_78;

	assign buf_78 = net_348;

	assign net_365 = buf_79;

	assign buf_79 = net_349;

	assign net_366 = buf_80;

	assign buf_80 = net_350;

	assign net_367 = buf_81;

	assign buf_81 = net_351;


	assign buf_82 = net_256;


	assign buf_83 = net_257;


	assign buf_84 = net_258;


	assign buf_85 = net_259;


	assign buf_86 = net_260;


	assign buf_87 = net_261;


	assign buf_88 = net_262;


	assign buf_89 = net_263;


	assign buf_90 = net_264;


	assign buf_91 = net_265;


	assign buf_92 = net_266;


	assign buf_93 = net_267;


	assign buf_94 = net_268;


	assign buf_95 = net_269;


	assign buf_96 = net_270;


	assign buf_97 = net_271;

	assign net_400 = buf_98;

	assign buf_98 = net_272;

	assign net_401 = buf_99;

	assign buf_99 = net_273;

	assign net_402 = buf_100;

	assign buf_100 = net_274;

	assign net_403 = buf_101;

	assign buf_101 = net_275;

	assign net_404 = buf_102;

	assign buf_102 = net_276;

	assign net_405 = buf_103;

	assign buf_103 = net_277;

	assign net_406 = buf_104;

	assign buf_104 = net_278;

	assign net_407 = buf_105;

	assign buf_105 = net_279;

	assign net_408 = buf_106;

	assign buf_106 = net_280;

	assign net_409 = buf_107;

	assign buf_107 = net_281;

	assign net_410 = buf_108;

	assign buf_108 = net_282;

	assign net_411 = buf_109;

	assign buf_109 = net_283;

	assign net_412 = buf_110;

	assign buf_110 = net_284;

	assign net_413 = buf_111;

	assign buf_111 = net_285;

	assign net_414 = buf_112;

	assign buf_112 = net_286;

	assign net_415 = buf_113;

	assign buf_113 = net_287;


	assign buf_114 = net_192;


	assign buf_115 = net_193;


	assign buf_116 = net_194;


	assign buf_117 = net_195;


	assign buf_118 = net_196;


	assign buf_119 = net_197;


	assign buf_120 = net_198;


	assign buf_121 = net_199;


	assign buf_122 = net_200;


	assign buf_123 = net_201;


	assign buf_124 = net_202;


	assign buf_125 = net_203;


	assign buf_126 = net_204;


	assign buf_127 = net_205;


	assign buf_128 = net_206;


	assign buf_129 = net_207;

	assign net_448 = buf_130;

	assign buf_130 = net_208;

	assign net_449 = buf_131;

	assign buf_131 = net_209;

	assign net_450 = buf_132;

	assign buf_132 = net_210;

	assign net_451 = buf_133;

	assign buf_133 = net_211;

	assign net_452 = buf_134;

	assign buf_134 = net_212;

	assign net_453 = buf_135;

	assign buf_135 = net_213;

	assign net_454 = buf_136;

	assign buf_136 = net_214;

	assign net_455 = buf_137;

	assign buf_137 = net_215;

	assign net_456 = buf_138;

	assign buf_138 = net_216;

	assign net_457 = buf_139;

	assign buf_139 = net_217;

	assign net_458 = buf_140;

	assign buf_140 = net_218;

	assign net_459 = buf_141;

	assign buf_141 = net_219;

	assign net_460 = buf_142;

	assign buf_142 = net_220;

	assign net_461 = buf_143;

	assign buf_143 = net_221;

	assign net_462 = buf_144;

	assign buf_144 = net_222;

	assign net_463 = buf_145;

	assign buf_145 = net_223;


	assign buf_146 = net_128;


	assign buf_147 = net_129;


	assign buf_148 = net_130;


	assign buf_149 = net_131;


	assign buf_150 = net_132;


	assign buf_151 = net_133;


	assign buf_152 = net_134;


	assign buf_153 = net_135;


	assign buf_154 = net_136;


	assign buf_155 = net_137;


	assign buf_156 = net_138;


	assign buf_157 = net_139;


	assign buf_158 = net_140;


	assign buf_159 = net_141;


	assign buf_160 = net_142;


	assign buf_161 = net_143;

	assign net_528 = buf_162;

	assign buf_162 = net_144;

	assign net_529 = buf_163;

	assign buf_163 = net_145;

	assign net_530 = buf_164;

	assign buf_164 = net_146;

	assign net_531 = buf_165;

	assign buf_165 = net_147;

	assign net_532 = buf_166;

	assign buf_166 = net_148;

	assign net_533 = buf_167;

	assign buf_167 = net_149;

	assign net_534 = buf_168;

	assign buf_168 = net_150;

	assign net_535 = buf_169;

	assign buf_169 = net_151;

	assign net_536 = buf_170;

	assign buf_170 = net_152;

	assign net_537 = buf_171;

	assign buf_171 = net_153;

	assign net_538 = buf_172;

	assign buf_172 = net_154;

	assign net_539 = buf_173;

	assign buf_173 = net_155;

	assign net_540 = buf_174;

	assign buf_174 = net_156;

	assign net_541 = buf_175;

	assign buf_175 = net_157;

	assign net_542 = buf_176;

	assign buf_176 = net_158;

	assign net_543 = buf_177;

	assign buf_177 = net_159;

	assign net_544 = buf_178;

	assign buf_178 = net_384;

	assign net_545 = buf_179;

	assign buf_179 = net_385;

	assign net_546 = buf_180;

	assign buf_180 = net_386;

	assign net_547 = buf_181;

	assign buf_181 = net_387;

	assign net_548 = buf_182;

	assign buf_182 = net_388;

	assign net_549 = buf_183;

	assign buf_183 = net_389;

	assign net_550 = buf_184;

	assign buf_184 = net_390;

	assign net_551 = buf_185;

	assign buf_185 = net_391;

	assign net_552 = buf_186;

	assign buf_186 = net_392;

	assign net_553 = buf_187;

	assign buf_187 = net_393;

	assign net_554 = buf_188;

	assign buf_188 = net_394;

	assign net_555 = buf_189;

	assign buf_189 = net_395;

	assign net_556 = buf_190;

	assign buf_190 = net_396;

	assign net_557 = buf_191;

	assign buf_191 = net_397;

	assign net_558 = buf_192;

	assign buf_192 = net_398;

	assign net_559 = buf_193;

	assign buf_193 = net_399;

	assign net_496 = buf_194;

	assign buf_194 = net_432;

	assign net_497 = buf_195;

	assign buf_195 = net_433;

	assign net_498 = buf_196;

	assign buf_196 = net_434;

	assign net_499 = buf_197;

	assign buf_197 = net_435;

	assign net_500 = buf_198;

	assign buf_198 = net_436;

	assign net_501 = buf_199;

	assign buf_199 = net_437;

	assign net_502 = buf_200;

	assign buf_200 = net_438;

	assign net_503 = buf_201;

	assign buf_201 = net_439;

	assign net_504 = buf_202;

	assign buf_202 = net_440;

	assign net_505 = buf_203;

	assign buf_203 = net_441;

	assign net_506 = buf_204;

	assign buf_204 = net_442;

	assign net_507 = buf_205;

	assign buf_205 = net_443;

	assign net_508 = buf_206;

	assign buf_206 = net_444;

	assign net_509 = buf_207;

	assign buf_207 = net_445;

	assign net_510 = buf_208;

	assign buf_208 = net_446;

	assign net_511 = buf_209;

	assign buf_209 = net_447;

	assign net_512 = buf_210;

	assign buf_210 = net_480;

	assign net_513 = buf_211;

	assign buf_211 = net_481;

	assign net_514 = buf_212;

	assign buf_212 = net_482;

	assign net_515 = buf_213;

	assign buf_213 = net_483;

	assign net_516 = buf_214;

	assign buf_214 = net_484;

	assign net_517 = buf_215;

	assign buf_215 = net_485;

	assign net_518 = buf_216;

	assign buf_216 = net_486;

	assign net_519 = buf_217;

	assign buf_217 = net_487;

	assign net_520 = buf_218;

	assign buf_218 = net_488;

	assign net_521 = buf_219;

	assign buf_219 = net_489;

	assign net_522 = buf_220;

	assign buf_220 = net_490;

	assign net_523 = buf_221;

	assign buf_221 = net_491;

	assign net_524 = buf_222;

	assign buf_222 = net_492;

	assign net_525 = buf_223;

	assign buf_223 = net_493;

	assign net_526 = buf_224;

	assign buf_224 = net_494;

	assign net_527 = buf_225;

	assign buf_225 = net_495;

	assign net_112 = buf_226;

	assign buf_226 = net_16;

	assign net_113 = buf_227;

	assign buf_227 = net_17;

	assign net_114 = buf_228;

	assign buf_228 = net_18;

	assign net_115 = buf_229;

	assign buf_229 = net_19;

	assign net_116 = buf_230;

	assign buf_230 = net_20;

	assign net_117 = buf_231;

	assign buf_231 = net_21;

	assign net_118 = buf_232;

	assign buf_232 = net_22;

	assign net_119 = buf_233;

	assign buf_233 = net_23;

	assign net_120 = buf_234;

	assign buf_234 = net_24;

	assign net_121 = buf_235;

	assign buf_235 = net_25;

	assign net_122 = buf_236;

	assign buf_236 = net_26;

	assign net_123 = buf_237;

	assign buf_237 = net_27;

	assign net_124 = buf_238;

	assign buf_238 = net_28;

	assign net_125 = buf_239;

	assign buf_239 = net_29;

	assign net_126 = buf_240;

	assign buf_240 = net_30;

	assign net_127 = buf_241;

	assign buf_241 = net_31;

	assign net_176 = buf_242;

	assign buf_242 = net_32;

	assign net_177 = buf_243;

	assign buf_243 = net_33;

	assign net_178 = buf_244;

	assign buf_244 = net_34;

	assign net_179 = buf_245;

	assign buf_245 = net_35;

	assign net_180 = buf_246;

	assign buf_246 = net_36;

	assign net_181 = buf_247;

	assign buf_247 = net_37;

	assign net_182 = buf_248;

	assign buf_248 = net_38;

	assign net_183 = buf_249;

	assign buf_249 = net_39;

	assign net_184 = buf_250;

	assign buf_250 = net_40;

	assign net_185 = buf_251;

	assign buf_251 = net_41;

	assign net_186 = buf_252;

	assign buf_252 = net_42;

	assign net_187 = buf_253;

	assign buf_253 = net_43;

	assign net_188 = buf_254;

	assign buf_254 = net_44;

	assign net_189 = buf_255;

	assign buf_255 = net_45;

	assign net_190 = buf_256;

	assign buf_256 = net_46;

	assign net_191 = buf_257;

	assign buf_257 = net_47;

	assign net_240 = buf_258;

	assign buf_258 = net_48;

	assign net_241 = buf_259;

	assign buf_259 = net_49;

	assign net_242 = buf_260;

	assign buf_260 = net_50;

	assign net_243 = buf_261;

	assign buf_261 = net_51;

	assign net_244 = buf_262;

	assign buf_262 = net_52;

	assign net_245 = buf_263;

	assign buf_263 = net_53;

	assign net_246 = buf_264;

	assign buf_264 = net_54;

	assign net_247 = buf_265;

	assign buf_265 = net_55;

	assign net_248 = buf_266;

	assign buf_266 = net_56;

	assign net_249 = buf_267;

	assign buf_267 = net_57;

	assign net_250 = buf_268;

	assign buf_268 = net_58;

	assign net_251 = buf_269;

	assign buf_269 = net_59;

	assign net_252 = buf_270;

	assign buf_270 = net_60;

	assign net_253 = buf_271;

	assign buf_271 = net_61;

	assign net_254 = buf_272;

	assign buf_272 = net_62;

	assign net_255 = buf_273;

	assign buf_273 = net_63;

	assign net_304 = buf_274;

	assign buf_274 = net_64;

	assign net_305 = buf_275;

	assign buf_275 = net_65;

	assign net_306 = buf_276;

	assign buf_276 = net_66;

	assign net_307 = buf_277;

	assign buf_277 = net_67;

	assign net_308 = buf_278;

	assign buf_278 = net_68;

	assign net_309 = buf_279;

	assign buf_279 = net_69;

	assign net_310 = buf_280;

	assign buf_280 = net_70;

	assign net_311 = buf_281;

	assign buf_281 = net_71;

	assign net_312 = buf_282;

	assign buf_282 = net_72;

	assign net_313 = buf_283;

	assign buf_283 = net_73;

	assign net_314 = buf_284;

	assign buf_284 = net_74;

	assign net_315 = buf_285;

	assign buf_285 = net_75;

	assign net_316 = buf_286;

	assign buf_286 = net_76;

	assign net_317 = buf_287;

	assign buf_287 = net_77;

	assign net_318 = buf_288;

	assign buf_288 = net_78;

	assign net_319 = buf_289;

	assign buf_289 = net_79;

	assign net_368 = q_290;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_290 = 1'b0;
		end
		else
		begin
			q_290 = net_496;
		end
	end

	assign net_369 = q_291;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_291 = 1'b0;
		end
		else
		begin
			q_291 = net_497;
		end
	end

	assign net_370 = q_292;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_292 = 1'b0;
		end
		else
		begin
			q_292 = net_498;
		end
	end

	assign net_371 = q_293;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_293 = 1'b0;
		end
		else
		begin
			q_293 = net_499;
		end
	end

	assign net_372 = q_294;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_294 = 1'b0;
		end
		else
		begin
			q_294 = net_500;
		end
	end

	assign net_373 = q_295;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_295 = 1'b0;
		end
		else
		begin
			q_295 = net_501;
		end
	end

	assign net_374 = q_296;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_296 = 1'b0;
		end
		else
		begin
			q_296 = net_502;
		end
	end

	assign net_375 = q_297;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_297 = 1'b0;
		end
		else
		begin
			q_297 = net_503;
		end
	end

	assign net_376 = q_298;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_298 = 1'b0;
		end
		else
		begin
			q_298 = net_504;
		end
	end

	assign net_377 = q_299;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_299 = 1'b0;
		end
		else
		begin
			q_299 = net_505;
		end
	end

	assign net_378 = q_300;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_300 = 1'b0;
		end
		else
		begin
			q_300 = net_506;
		end
	end

	assign net_379 = q_301;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_301 = 1'b0;
		end
		else
		begin
			q_301 = net_507;
		end
	end

	assign net_380 = q_302;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_302 = 1'b0;
		end
		else
		begin
			q_302 = net_508;
		end
	end

	assign net_381 = q_303;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_303 = 1'b0;
		end
		else
		begin
			q_303 = net_509;
		end
	end

	assign net_382 = q_304;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_304 = 1'b0;
		end
		else
		begin
			q_304 = net_510;
		end
	end

	assign net_383 = q_305;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_305 = 1'b0;
		end
		else
		begin
			q_305 = net_511;
		end
	end

	assign net_416 = q_306;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_306 = 1'b0;
		end
		else
		begin
			q_306 = net_512;
		end
	end

	assign net_417 = q_307;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_307 = 1'b0;
		end
		else
		begin
			q_307 = net_513;
		end
	end

	assign net_418 = q_308;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_308 = 1'b0;
		end
		else
		begin
			q_308 = net_514;
		end
	end

	assign net_419 = q_309;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_309 = 1'b0;
		end
		else
		begin
			q_309 = net_515;
		end
	end

	assign net_420 = q_310;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_310 = 1'b0;
		end
		else
		begin
			q_310 = net_516;
		end
	end

	assign net_421 = q_311;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_311 = 1'b0;
		end
		else
		begin
			q_311 = net_517;
		end
	end

	assign net_422 = q_312;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_312 = 1'b0;
		end
		else
		begin
			q_312 = net_518;
		end
	end

	assign net_423 = q_313;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_313 = 1'b0;
		end
		else
		begin
			q_313 = net_519;
		end
	end

	assign net_424 = q_314;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_314 = 1'b0;
		end
		else
		begin
			q_314 = net_520;
		end
	end

	assign net_425 = q_315;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_315 = 1'b0;
		end
		else
		begin
			q_315 = net_521;
		end
	end

	assign net_426 = q_316;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_316 = 1'b0;
		end
		else
		begin
			q_316 = net_522;
		end
	end

	assign net_427 = q_317;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_317 = 1'b0;
		end
		else
		begin
			q_317 = net_523;
		end
	end

	assign net_428 = q_318;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_318 = 1'b0;
		end
		else
		begin
			q_318 = net_524;
		end
	end

	assign net_429 = q_319;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_319 = 1'b0;
		end
		else
		begin
			q_319 = net_525;
		end
	end

	assign net_430 = q_320;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_320 = 1'b0;
		end
		else
		begin
			q_320 = net_526;
		end
	end

	assign net_431 = q_321;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_321 = 1'b0;
		end
		else
		begin
			q_321 = net_527;
		end
	end

	assign net_464 = q_322;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_322 = 1'b0;
		end
		else
		begin
			q_322 = net_528;
		end
	end

	assign net_465 = q_323;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_323 = 1'b0;
		end
		else
		begin
			q_323 = net_529;
		end
	end

	assign net_466 = q_324;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_324 = 1'b0;
		end
		else
		begin
			q_324 = net_530;
		end
	end

	assign net_467 = q_325;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_325 = 1'b0;
		end
		else
		begin
			q_325 = net_531;
		end
	end

	assign net_468 = q_326;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_326 = 1'b0;
		end
		else
		begin
			q_326 = net_532;
		end
	end

	assign net_469 = q_327;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_327 = 1'b0;
		end
		else
		begin
			q_327 = net_533;
		end
	end

	assign net_470 = q_328;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_328 = 1'b0;
		end
		else
		begin
			q_328 = net_534;
		end
	end

	assign net_471 = q_329;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_329 = 1'b0;
		end
		else
		begin
			q_329 = net_535;
		end
	end

	assign net_472 = q_330;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_330 = 1'b0;
		end
		else
		begin
			q_330 = net_536;
		end
	end

	assign net_473 = q_331;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_331 = 1'b0;
		end
		else
		begin
			q_331 = net_537;
		end
	end

	assign net_474 = q_332;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_332 = 1'b0;
		end
		else
		begin
			q_332 = net_538;
		end
	end

	assign net_475 = q_333;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_333 = 1'b0;
		end
		else
		begin
			q_333 = net_539;
		end
	end

	assign net_476 = q_334;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_334 = 1'b0;
		end
		else
		begin
			q_334 = net_540;
		end
	end

	assign net_477 = q_335;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_335 = 1'b0;
		end
		else
		begin
			q_335 = net_541;
		end
	end

	assign net_478 = q_336;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_336 = 1'b0;
		end
		else
		begin
			q_336 = net_542;
		end
	end

	assign net_479 = q_337;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_337 = 1'b0;
		end
		else
		begin
			q_337 = net_543;
		end
	end

	assign net_96 = q_338;
	assign net_160 = q_338;
	assign net_224 = q_338;
	assign net_288 = q_338;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_338 = 1'b0;
		end
		else
		begin
			q_338 = net_80;
		end
	end

	assign net_97 = q_339;
	assign net_161 = q_339;
	assign net_225 = q_339;
	assign net_289 = q_339;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_339 = 1'b0;
		end
		else
		begin
			q_339 = net_81;
		end
	end

	assign net_98 = q_340;
	assign net_162 = q_340;
	assign net_226 = q_340;
	assign net_290 = q_340;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_340 = 1'b0;
		end
		else
		begin
			q_340 = net_82;
		end
	end

	assign net_99 = q_341;
	assign net_163 = q_341;
	assign net_227 = q_341;
	assign net_291 = q_341;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_341 = 1'b0;
		end
		else
		begin
			q_341 = net_83;
		end
	end

	assign net_100 = q_342;
	assign net_164 = q_342;
	assign net_228 = q_342;
	assign net_292 = q_342;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_342 = 1'b0;
		end
		else
		begin
			q_342 = net_84;
		end
	end

	assign net_101 = q_343;
	assign net_165 = q_343;
	assign net_229 = q_343;
	assign net_293 = q_343;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_343 = 1'b0;
		end
		else
		begin
			q_343 = net_85;
		end
	end

	assign net_102 = q_344;
	assign net_166 = q_344;
	assign net_230 = q_344;
	assign net_294 = q_344;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_344 = 1'b0;
		end
		else
		begin
			q_344 = net_86;
		end
	end

	assign net_103 = q_345;
	assign net_167 = q_345;
	assign net_231 = q_345;
	assign net_295 = q_345;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_345 = 1'b0;
		end
		else
		begin
			q_345 = net_87;
		end
	end

	assign net_104 = q_346;
	assign net_168 = q_346;
	assign net_232 = q_346;
	assign net_296 = q_346;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_346 = 1'b0;
		end
		else
		begin
			q_346 = net_88;
		end
	end

	assign net_105 = q_347;
	assign net_169 = q_347;
	assign net_233 = q_347;
	assign net_297 = q_347;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_347 = 1'b0;
		end
		else
		begin
			q_347 = net_89;
		end
	end

	assign net_106 = q_348;
	assign net_170 = q_348;
	assign net_234 = q_348;
	assign net_298 = q_348;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_348 = 1'b0;
		end
		else
		begin
			q_348 = net_90;
		end
	end

	assign net_107 = q_349;
	assign net_171 = q_349;
	assign net_235 = q_349;
	assign net_299 = q_349;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_349 = 1'b0;
		end
		else
		begin
			q_349 = net_91;
		end
	end

	assign net_108 = q_350;
	assign net_172 = q_350;
	assign net_236 = q_350;
	assign net_300 = q_350;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_350 = 1'b0;
		end
		else
		begin
			q_350 = net_92;
		end
	end

	assign net_109 = q_351;
	assign net_173 = q_351;
	assign net_237 = q_351;
	assign net_301 = q_351;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_351 = 1'b0;
		end
		else
		begin
			q_351 = net_93;
		end
	end

	assign net_110 = q_352;
	assign net_174 = q_352;
	assign net_238 = q_352;
	assign net_302 = q_352;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_352 = 1'b0;
		end
		else
		begin
			q_352 = net_94;
		end
	end

	assign net_111 = q_353;
	assign net_175 = q_353;
	assign net_239 = q_353;
	assign net_303 = q_353;

	always@(posedge clk, posedge rst)
	begin
		if (rst)
		begin
			q_353 = 1'b0;
		end
		else
		begin
			q_353 = net_95;
		end
	end

	assign net_128 = mult_354[0];
	assign net_129 = mult_354[1];
	assign net_130 = mult_354[2];
	assign net_131 = mult_354[3];
	assign net_132 = mult_354[4];
	assign net_133 = mult_354[5];
	assign net_134 = mult_354[6];
	assign net_135 = mult_354[7];
	assign net_136 = mult_354[8];
	assign net_137 = mult_354[9];
	assign net_138 = mult_354[10];
	assign net_139 = mult_354[11];
	assign net_140 = mult_354[12];
	assign net_141 = mult_354[13];
	assign net_142 = mult_354[14];
	assign net_143 = mult_354[15];
	assign net_144 = mult_354[16];
	assign net_145 = mult_354[17];
	assign net_146 = mult_354[18];
	assign net_147 = mult_354[19];
	assign net_148 = mult_354[20];
	assign net_149 = mult_354[21];
	assign net_150 = mult_354[22];
	assign net_151 = mult_354[23];
	assign net_152 = mult_354[24];
	assign net_153 = mult_354[25];
	assign net_154 = mult_354[26];
	assign net_155 = mult_354[27];
	assign net_156 = mult_354[28];
	assign net_157 = mult_354[29];
	assign net_158 = mult_354[30];
	assign net_159 = mult_354[31];

	assign mult_354 = {net_111, net_110, net_109, net_108, net_107, net_106, net_105, net_104, net_103, net_102, net_101, net_100, net_99, net_98, net_97, net_96} * {net_127, net_126, net_125, net_124, net_123, net_122, net_121, net_120, net_119, net_118, net_117, net_116, net_115, net_114, net_113, net_112};

	assign net_192 = mult_355[0];
	assign net_193 = mult_355[1];
	assign net_194 = mult_355[2];
	assign net_195 = mult_355[3];
	assign net_196 = mult_355[4];
	assign net_197 = mult_355[5];
	assign net_198 = mult_355[6];
	assign net_199 = mult_355[7];
	assign net_200 = mult_355[8];
	assign net_201 = mult_355[9];
	assign net_202 = mult_355[10];
	assign net_203 = mult_355[11];
	assign net_204 = mult_355[12];
	assign net_205 = mult_355[13];
	assign net_206 = mult_355[14];
	assign net_207 = mult_355[15];
	assign net_208 = mult_355[16];
	assign net_209 = mult_355[17];
	assign net_210 = mult_355[18];
	assign net_211 = mult_355[19];
	assign net_212 = mult_355[20];
	assign net_213 = mult_355[21];
	assign net_214 = mult_355[22];
	assign net_215 = mult_355[23];
	assign net_216 = mult_355[24];
	assign net_217 = mult_355[25];
	assign net_218 = mult_355[26];
	assign net_219 = mult_355[27];
	assign net_220 = mult_355[28];
	assign net_221 = mult_355[29];
	assign net_222 = mult_355[30];
	assign net_223 = mult_355[31];

	assign mult_355 = {net_175, net_174, net_173, net_172, net_171, net_170, net_169, net_168, net_167, net_166, net_165, net_164, net_163, net_162, net_161, net_160} * {net_191, net_190, net_189, net_188, net_187, net_186, net_185, net_184, net_183, net_182, net_181, net_180, net_179, net_178, net_177, net_176};

	assign net_256 = mult_356[0];
	assign net_257 = mult_356[1];
	assign net_258 = mult_356[2];
	assign net_259 = mult_356[3];
	assign net_260 = mult_356[4];
	assign net_261 = mult_356[5];
	assign net_262 = mult_356[6];
	assign net_263 = mult_356[7];
	assign net_264 = mult_356[8];
	assign net_265 = mult_356[9];
	assign net_266 = mult_356[10];
	assign net_267 = mult_356[11];
	assign net_268 = mult_356[12];
	assign net_269 = mult_356[13];
	assign net_270 = mult_356[14];
	assign net_271 = mult_356[15];
	assign net_272 = mult_356[16];
	assign net_273 = mult_356[17];
	assign net_274 = mult_356[18];
	assign net_275 = mult_356[19];
	assign net_276 = mult_356[20];
	assign net_277 = mult_356[21];
	assign net_278 = mult_356[22];
	assign net_279 = mult_356[23];
	assign net_280 = mult_356[24];
	assign net_281 = mult_356[25];
	assign net_282 = mult_356[26];
	assign net_283 = mult_356[27];
	assign net_284 = mult_356[28];
	assign net_285 = mult_356[29];
	assign net_286 = mult_356[30];
	assign net_287 = mult_356[31];

	assign mult_356 = {net_239, net_238, net_237, net_236, net_235, net_234, net_233, net_232, net_231, net_230, net_229, net_228, net_227, net_226, net_225, net_224} * {net_255, net_254, net_253, net_252, net_251, net_250, net_249, net_248, net_247, net_246, net_245, net_244, net_243, net_242, net_241, net_240};

	assign net_320 = mult_357[0];
	assign net_321 = mult_357[1];
	assign net_322 = mult_357[2];
	assign net_323 = mult_357[3];
	assign net_324 = mult_357[4];
	assign net_325 = mult_357[5];
	assign net_326 = mult_357[6];
	assign net_327 = mult_357[7];
	assign net_328 = mult_357[8];
	assign net_329 = mult_357[9];
	assign net_330 = mult_357[10];
	assign net_331 = mult_357[11];
	assign net_332 = mult_357[12];
	assign net_333 = mult_357[13];
	assign net_334 = mult_357[14];
	assign net_335 = mult_357[15];
	assign net_336 = mult_357[16];
	assign net_337 = mult_357[17];
	assign net_338 = mult_357[18];
	assign net_339 = mult_357[19];
	assign net_340 = mult_357[20];
	assign net_341 = mult_357[21];
	assign net_342 = mult_357[22];
	assign net_343 = mult_357[23];
	assign net_344 = mult_357[24];
	assign net_345 = mult_357[25];
	assign net_346 = mult_357[26];
	assign net_347 = mult_357[27];
	assign net_348 = mult_357[28];
	assign net_349 = mult_357[29];
	assign net_350 = mult_357[30];
	assign net_351 = mult_357[31];

	assign mult_357 = {net_303, net_302, net_301, net_300, net_299, net_298, net_297, net_296, net_295, net_294, net_293, net_292, net_291, net_290, net_289, net_288} * {net_319, net_318, net_317, net_316, net_315, net_314, net_313, net_312, net_311, net_310, net_309, net_308, net_307, net_306, net_305, net_304};

	assign net_384 = add_358[0];
	assign net_385 = add_358[1];
	assign net_386 = add_358[2];
	assign net_387 = add_358[3];
	assign net_388 = add_358[4];
	assign net_389 = add_358[5];
	assign net_390 = add_358[6];
	assign net_391 = add_358[7];
	assign net_392 = add_358[8];
	assign net_393 = add_358[9];
	assign net_394 = add_358[10];
	assign net_395 = add_358[11];
	assign net_396 = add_358[12];
	assign net_397 = add_358[13];
	assign net_398 = add_358[14];
	assign net_399 = add_358[15];

	assign add_358 = {net_367, net_366, net_365, net_364, net_363, net_362, net_361, net_360, net_359, net_358, net_357, net_356, net_355, net_354, net_353, net_352} + {net_383, net_382, net_381, net_380, net_379, net_378, net_377, net_376, net_375, net_374, net_373, net_372, net_371, net_370, net_369, net_368};

	assign net_432 = add_359[0];
	assign net_433 = add_359[1];
	assign net_434 = add_359[2];
	assign net_435 = add_359[3];
	assign net_436 = add_359[4];
	assign net_437 = add_359[5];
	assign net_438 = add_359[6];
	assign net_439 = add_359[7];
	assign net_440 = add_359[8];
	assign net_441 = add_359[9];
	assign net_442 = add_359[10];
	assign net_443 = add_359[11];
	assign net_444 = add_359[12];
	assign net_445 = add_359[13];
	assign net_446 = add_359[14];
	assign net_447 = add_359[15];

	assign add_359 = {net_415, net_414, net_413, net_412, net_411, net_410, net_409, net_408, net_407, net_406, net_405, net_404, net_403, net_402, net_401, net_400} + {net_431, net_430, net_429, net_428, net_427, net_426, net_425, net_424, net_423, net_422, net_421, net_420, net_419, net_418, net_417, net_416};

	assign net_480 = add_360[0];
	assign net_481 = add_360[1];
	assign net_482 = add_360[2];
	assign net_483 = add_360[3];
	assign net_484 = add_360[4];
	assign net_485 = add_360[5];
	assign net_486 = add_360[6];
	assign net_487 = add_360[7];
	assign net_488 = add_360[8];
	assign net_489 = add_360[9];
	assign net_490 = add_360[10];
	assign net_491 = add_360[11];
	assign net_492 = add_360[12];
	assign net_493 = add_360[13];
	assign net_494 = add_360[14];
	assign net_495 = add_360[15];

	assign add_360 = {net_463, net_462, net_461, net_460, net_459, net_458, net_457, net_456, net_455, net_454, net_453, net_452, net_451, net_450, net_449, net_448} + {net_479, net_478, net_477, net_476, net_475, net_474, net_473, net_472, net_471, net_470, net_469, net_468, net_467, net_466, net_465, net_464};

endmodule
